* Title: Test circuit

* Netlist
R0 n22 0 0
D3 n22 n21 DMOD
.model DMOD D
R4 n25 n21 470000.0
D6 n21 n22 DMOD
.model DMOD D
C10 n25 n27 0.22 ic=0.0
R13 n27 n25 160.0
V14 n27 n28 SIN(0.0 230.0 50.0 0.001 0.0 0.0)
R15 n28 0 0

.control
op
tran 0.1 0.2 0 uic
echo output test > result.txt $ start new file
set appendwrite
set wr_vecnames
set wr_singlescale
wrdata data.txt all
.endc
