* Title: Test circuit

* Netlist
R1 n18 0 0
R3 n20 n21 470000.0
D4 n18 n21 DMOD
.model DMOD D
D7 n21 n18 DMOD
.model DMOD D
C10 n20 n26 0.22 ic=0.0
R13 n26 n20 160.0
V14 n26 n28 SIN(0.0 230.0 50.0 0.001 0.0 0.0)
R15 n28 0 0

.control
op
tran 1.0 0.4 0 uic
echo output test > result.txt $ start new file
set appendwrite
set wr_vecnames
set wr_singlescale
wrdata data.txt all
.endc
