* Title: Test circuit

* Netlist
V0 n32 n26 5.0
D3 n25 n19 DMOD
.model DMOD D
Q4 n33 n19 n29 QMOD
.model QMOD NPN level=4
R7 n29 0 0
R10 n24 0 0
V11 n19 n24 SIN(0.0 1.0 0.0 0.001 0.0 0.0)
R12 n25 0 0
R13 n26 0 0
R17 n32 n33 10.0

.control
op
tran 0.1 5.0 0 uic
echo output test > result.txt $ start new file
set appendwrite
set wr_vecnames
set wr_singlescale
wrdata data.txt all
.endc
