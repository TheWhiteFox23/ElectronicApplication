* Title: Test circuit

* Netlist
V1 n25 n19 5.0
Q2 n22 n21 n26 QMOD
.model QMOD PNP level=4
R5 n22 0 0
R7 n18 0 0
V8 n21 n18 SIN(0.0 1.0 0.0 0.001 0.0 0.0)
R9 n19 0 0
R13 n25 n26 10.0

.control
op
tran 0.1 5.0 0 uic
echo output test > result.txt $ start new file
set appendwrite
set wr_vecnames
set wr_singlescale
wrdata data.txt all
.endc
